module Shifter( result, leftRight, shamt, sftSrc );

//I/O ports 
input	leftRight;
input	[32-1:0] shamt;
input	[32-1:0] sftSrc ;

output	[32-1:0] result;
//Internal Signals
wire	[32-1:0] result;
  
//Main function
/*your code here*/

assign result = 	(!leftRight)?(sftSrc>>shamt):	//rightshift if 0
						(leftRight)?(sftSrc<<shamt):
						32'd0;//default

endmodule